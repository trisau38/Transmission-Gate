magic
tech scmos
timestamp 1664282788
<< nwell >>
rect -19 -5 6 31
<< polysilicon >>
rect -9 21 -5 33
rect -9 -5 -5 -3
rect -9 -14 -5 -11
rect -9 -25 -5 -22
<< ndiffusion >>
rect -17 -16 -9 -14
rect -17 -20 -15 -16
rect -11 -20 -9 -16
rect -17 -22 -9 -20
rect -5 -16 4 -14
rect -5 -20 -2 -16
rect 2 -20 4 -16
rect -5 -22 4 -20
<< pdiffusion >>
rect -17 11 -9 21
rect -17 7 -15 11
rect -11 7 -9 11
rect -17 -3 -9 7
rect -5 11 4 21
rect -5 7 -2 11
rect 2 7 4 11
rect -5 -3 4 7
<< metal1 >>
rect -35 40 24 44
rect -9 37 -5 40
rect 3 25 15 29
rect -15 -16 -11 7
rect -9 -32 -5 -29
rect 11 -32 15 25
rect -35 -36 24 -32
<< metal2 >>
rect -2 -20 2 11
<< ntransistor >>
rect -9 -22 -5 -14
<< ptransistor >>
rect -9 -3 -5 21
<< polycontact >>
rect -9 33 -5 37
rect -9 -29 -5 -25
<< ndcontact >>
rect -15 -20 -11 -16
rect -2 -20 2 -16
<< pdcontact >>
rect -15 7 -11 11
rect -2 7 2 11
<< nsubstratencontact >>
rect -1 25 3 29
<< labels >>
rlabel metal1 -7 -34 -7 -34 1 VDD
rlabel metal1 -13 -10 -13 -10 1 in
rlabel metal2 0 -9 0 -9 1 out
rlabel metal1 -7 42 -7 42 5 GND
<< end >>
